// Author: Dylan Boland
//
// Parameters used throughout the design.

parameter TRFC_PB_WIDTH = 4;
parameter BANK_ADDR_WIDTH = 4;