// Author: Dylan Boland
//
//
`include "design_parameters.svh" // include the design parameters

module tRFCpb_checker #
	(
	// ==== Parameters ====
	parameter NUM_TRFC_PB_CNTRS = 4,
	parameter NUM_BANKS = 16
	)
	(
	// ==== Inputs ====
	input logic clk,
	input logic rst_n,
	input logic refpb_issued,
	// ==== Outputs ====
	output logic [NUM_BANKS-1:0] trfc_pb_met // indicates which banks have met the tRFCpb time requirement
	);

	// ==== Signal Declarations ====
	logic [NUM_TRFC_PB_CNTRS-1:0] trfc_pb_cntrs_assigned;
	// The signal below will be generated by inverting each bit
	// in the signal above (trfc_pb_cntrs_assigned):
	logic [NUM_TRFC_PB_CNTRS-1:0] trfc_pb_cntrs_available;
	logic trfc_pb_cntr_free; // generated by OR-ing all the bits in trfc_pb_cntrs_available
	logic [NUM_TRFC_PB_CNTRS-1:0] trfc_pb_cntrs_elapsed;
	logic trfc_pb_cntr_elapsed; // equal to the OR of all the bits in trfc_pb_cntrs_elapsed
	logic [NUM_BANKS-1:0] trfc_pb_met; // indicates which banks have met the tRFCpb time requirement
	logic [NUM_TRFC_PB_CNTRS-1:0] trfc_pb_cntr_triggers;
	logic [NUM_BANKS-1:0] banks_available_for_refresh; // indicates which banks can be refreshed
	// The signal below indicates which counter has been selected to
	// measure the tRFCpb time. For example, if there were two counters, and
	// the signal were equal to 2'b01, it would indicate that the first counter
	// was selected to measure the tRFCpb time. If the signal were set to 2'b10
	// then it would indicate that the second counter was chosen. Importantly, only
	// one bit will be set in this signal.
	logic [NUM_TRFC_PB_CNTRS-1:0] selected_trfc_pb_cntr;
	// The signal below has "NUM_TRFC_PB_CNTRS" segments, with each segments
	// having a width equal to "BANK_ADDR_WIDTH". It indicates which bank (if any)
	// is assigned to each tRFCpb counter (timer):
	logic [NUM_TRFC_PB_CNTRS-1:0][BANK_ADDR_WIDTH-1:0] bank_assigned_trfc_pb_cntr;
	// The bus signal below is driven by the tRFCpb counters.
	logic [NUM_TRFC_PB_CNTRS-1:0][BANK_ADDR_WIDTH-1:0] assigned_bank_trfc_pb_cntr;

	// ==== Signal Definitions ====
	assign trfc_pb_cntrs_available = ~trfc_pb_cntrs_assigned;
	assign trfc_pb_cntr_elapsed = |trfc_pb_cntrs_elapsed;

	// ==== Logic for choosing which counter will be used ====
	always_comb begin
		selected_trfc_pb_cntr = {NUM_TRFC_PB_CNTRS{1'b0}};
		for (int i = 0; i < NUM_TRFC_PB_CNTRS; i = i + 1) begin
			if (trfc_pb_cntrs_available[i]) begin
				selected_trfc_pb_cntr[i] = 1'b1;
				break;
			end
		end
	end

	// ==== Logic for generating the counter-trigger signals (i.e., start signals) ====
	assign trfc_pb_cntr_triggers = selected_trfc_pb_cntr & {NUM_TRFC_PB_CNTRS{refpb_issued}};

	// ==== Instantiate the Refresh-Cycle-Time (tRFCpb) Counters ====
	genvar n;
	generate
		for (n = 0; n < NUM_TRFC_PB_CNTRS; n = n + 1) begin: instantiate_tRFCpb_counters
			refresh_cycle_time_counter tRFCpb_timer
			(
			// ==== Inputs ====
			.clk(clk),
			.rst_n(rst_n),
			.start(trfc_pb_cntr_triggers[n]), // route the relevant bit of the "trigger" bus to the "start" input
			.trfc_pb(trfc_pb),
			.bank_assigned(bank_assigned_trfc_pb_cntr[n]), // route the right part of the bank_assigned_trfc_pb_cntr bus into the bank_assigned port
			// ==== Outputs ====
			.assigned(trfc_pb_cntrs_assigned[n]),
			.counter_done(trfc_pb_cntrs_elapsed[n]),
			.assigned_bank(assigned_bank_trfc_pb_cntr[n])
			);
		end
	endgenerate

endmodule






